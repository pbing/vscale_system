/* POCI type definitions */

package pk_poci;
   parameter
     data_width = 32,
     addr_width = 32;
endpackage
